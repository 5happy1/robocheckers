module not_32(in, out);

input [31:0] in;
output [31:0] out;

not not_0(out[0], in[0]);
not not_1(out[1], in[1]);
not not_2(out[2], in[2]);
not not_3(out[3], in[3]);
not not_4(out[4], in[4]);
not not_5(out[5], in[5]);
not not_6(out[6], in[6]);
not not_7(out[7], in[7]);
not not_8(out[8], in[8]);
not not_9(out[9], in[9]);
not not_10(out[10], in[10]);
not not_11(out[11], in[11]);
not not_12(out[12], in[12]);
not not_13(out[13], in[13]);
not not_14(out[14], in[14]);
not not_15(out[15], in[15]);
not not_16(out[16], in[16]);
not not_17(out[17], in[17]);
not not_18(out[18], in[18]);
not not_19(out[19], in[19]);
not not_20(out[20], in[20]);
not not_21(out[21], in[21]);
not not_22(out[22], in[22]);
not not_23(out[23], in[23]);
not not_24(out[24], in[24]);
not not_25(out[25], in[25]);
not not_26(out[26], in[26]);
not not_27(out[27], in[27]);
not not_28(out[28], in[28]);
not not_29(out[29], in[29]);
not not_30(out[30], in[30]);
not not_31(out[31], in[31]);

endmodule
