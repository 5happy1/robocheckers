module test_serial(data_in, data_out, clock_out);

input data_in, clock_in;
output data_out, clock_out;

derial d0(data_in, clock_in, data_out, clock_out);



endmodule
