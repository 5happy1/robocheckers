module and_32(in1, in2, out);

input [31:0] in1, in2;
output [31:0] out;

and and_0(out[0], in1[0], in2[0]);
and and_1(out[1], in1[1], in2[1]);
and and_2(out[2], in1[2], in2[2]);
and and_3(out[3], in1[3], in2[3]);
and and_4(out[4], in1[4], in2[4]);
and and_5(out[5], in1[5], in2[5]);
and and_6(out[6], in1[6], in2[6]);
and and_7(out[7], in1[7], in2[7]);
and and_8(out[8], in1[8], in2[8]);
and and_9(out[9], in1[9], in2[9]);
and and_10(out[10], in1[10], in2[10]);
and and_11(out[11], in1[11], in2[11]);
and and_12(out[12], in1[12], in2[12]);
and and_13(out[13], in1[13], in2[13]);
and and_14(out[14], in1[14], in2[14]);
and and_15(out[15], in1[15], in2[15]);
and and_16(out[16], in1[16], in2[16]);
and and_17(out[17], in1[17], in2[17]);
and and_18(out[18], in1[18], in2[18]);
and and_19(out[19], in1[19], in2[19]);
and and_20(out[20], in1[20], in2[20]);
and and_21(out[21], in1[21], in2[21]);
and and_22(out[22], in1[22], in2[22]);
and and_23(out[23], in1[23], in2[23]);
and and_24(out[24], in1[24], in2[24]);
and and_25(out[25], in1[25], in2[25]);
and and_26(out[26], in1[26], in2[26]);
and and_27(out[27], in1[27], in2[27]);
and and_28(out[28], in1[28], in2[28]);
and and_29(out[29], in1[29], in2[29]);
and and_30(out[30], in1[30], in2[30]);
and and_31(out[31], in1[31], in2[31]);

endmodule
