module mux_32(in, select, out);

input [31:0] in;
input [4:0] select;
output out;

endmodule
