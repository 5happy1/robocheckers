module comp_32(in1, in2, eq_out, gt_out);

input [31:0] in1, in2;
output eq_out, gt_out;

wire eq_15, gt_15;
wire eq_14, gt_14;
wire eq_13, gt_13;
wire eq_12, gt_12;
wire eq_11, gt_11;
wire eq_10, gt_10;
wire eq_9, gt_9;
wire eq_8, gt_8;
wire eq_7, gt_7;
wire eq_6, gt_6;
wire eq_5, gt_5;
wire eq_4, gt_4;
wire eq_3, gt_3;
wire eq_2, gt_2;
wire eq_1, gt_1;
wire eq_0, gt_0;

//comp_2 comp_15(eq_15

endmodule
